-- $Header: $
-------------------------------------------------------
--  Copyright (c) 2011 Xilinx Inc.
--  All Right Reserved.
-------------------------------------------------------
--
--   ____  ____
--  /   /\/   / 
-- /___/  \  /     Vendor      : Xilinx 
-- \   \   \/      Version     : 2012.2 
--  \   \          Description : 
--  /   /                      
-- /___/   /\      Filename    : MUXF9.vhd
-- \   \  /  \      
--  \__ \/\__ \                   
--                                 
--  Generated by    : /home/unified/chen/g2ltw/g2ltw.pl
--  Revision: 1.0
-------------------------------------------------------

----- CELL MUXF9 -----

library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity MUXF9 is
  port (
    O                    : out std_ulogic;
    I0                   : in std_ulogic;
    I1                   : in std_ulogic;
    S                    : in std_ulogic      
  );
end MUXF9;

architecture MUXF9_V of MUXF9 is
begin
  FunctionalBehavior   : process (I0, I1, S)
  begin
    if (S = '0') then
      O <= I0;
    else
      O <= I1;
    end if;
  end process;
end MUXF9_V;
