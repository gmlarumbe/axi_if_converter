-- $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/vhdsclibs/data/unisims/pele/VITAL/PS7.vhd,v 1.3 2011/04/28 18:02:53 harikr Exp $
-------------------------------------------------------
--  Copyright (c) 2011 Xilinx Inc.
--  All Right Reserved.
-------------------------------------------------------
--
--   ____  ____
--  /   /\/   / 
-- /___/  \  /     Vendor      : Xilinx 
-- \   \   \/      Version     : 13.1 
--  \   \          Description : 
--  /   /                      
-- /___/   /\      Filename    : PS7.vhd
-- \   \  /  \      
--  \__ \/\__ \                   
--                                 
--  Generated by    : /home/chen/xfoundry/HEAD/env/Databases/CAEInterfaces/LibraryWriters/bin/ltw.pl
--  Revision: 1.0
--  05/13/13 - 717829 - Add simulation message
-------------------------------------------------------

----- CELL PS7 -----

library IEEE;
use IEEE.STD_LOGIC_arith.all;
use IEEE.STD_LOGIC_1164.all;

library STD;
use STD.TEXTIO.all;

library unisim;
use unisim.VCOMPONENTS.all;
use unisim.vpkg.all;

  entity PS7 is
    port (
      DMA0DATYPE           : out std_logic_vector(1 downto 0);
      DMA0DAVALID          : out std_ulogic;
      DMA0DRREADY          : out std_ulogic;
      DMA0RSTN             : out std_ulogic;
      DMA1DATYPE           : out std_logic_vector(1 downto 0);
      DMA1DAVALID          : out std_ulogic;
      DMA1DRREADY          : out std_ulogic;
      DMA1RSTN             : out std_ulogic;
      DMA2DATYPE           : out std_logic_vector(1 downto 0);
      DMA2DAVALID          : out std_ulogic;
      DMA2DRREADY          : out std_ulogic;
      DMA2RSTN             : out std_ulogic;
      DMA3DATYPE           : out std_logic_vector(1 downto 0);
      DMA3DAVALID          : out std_ulogic;
      DMA3DRREADY          : out std_ulogic;
      DMA3RSTN             : out std_ulogic;
      EMIOCAN0PHYTX        : out std_ulogic;
      EMIOCAN1PHYTX        : out std_ulogic;
      EMIOENET0GMIITXD     : out std_logic_vector(7 downto 0);
      EMIOENET0GMIITXEN    : out std_ulogic;
      EMIOENET0GMIITXER    : out std_ulogic;
      EMIOENET0MDIOMDC     : out std_ulogic;
      EMIOENET0MDIOO       : out std_ulogic;
      EMIOENET0MDIOTN      : out std_ulogic;
      EMIOENET0PTPDELAYREQRX : out std_ulogic;
      EMIOENET0PTPDELAYREQTX : out std_ulogic;
      EMIOENET0PTPPDELAYREQRX : out std_ulogic;
      EMIOENET0PTPPDELAYREQTX : out std_ulogic;
      EMIOENET0PTPPDELAYRESPRX : out std_ulogic;
      EMIOENET0PTPPDELAYRESPTX : out std_ulogic;
      EMIOENET0PTPSYNCFRAMERX : out std_ulogic;
      EMIOENET0PTPSYNCFRAMETX : out std_ulogic;
      EMIOENET0SOFRX       : out std_ulogic;
      EMIOENET0SOFTX       : out std_ulogic;
      EMIOENET1GMIITXD     : out std_logic_vector(7 downto 0);
      EMIOENET1GMIITXEN    : out std_ulogic;
      EMIOENET1GMIITXER    : out std_ulogic;
      EMIOENET1MDIOMDC     : out std_ulogic;
      EMIOENET1MDIOO       : out std_ulogic;
      EMIOENET1MDIOTN      : out std_ulogic;
      EMIOENET1PTPDELAYREQRX : out std_ulogic;
      EMIOENET1PTPDELAYREQTX : out std_ulogic;
      EMIOENET1PTPPDELAYREQRX : out std_ulogic;
      EMIOENET1PTPPDELAYREQTX : out std_ulogic;
      EMIOENET1PTPPDELAYRESPRX : out std_ulogic;
      EMIOENET1PTPPDELAYRESPTX : out std_ulogic;
      EMIOENET1PTPSYNCFRAMERX : out std_ulogic;
      EMIOENET1PTPSYNCFRAMETX : out std_ulogic;
      EMIOENET1SOFRX       : out std_ulogic;
      EMIOENET1SOFTX       : out std_ulogic;
      EMIOGPIOO            : out std_logic_vector(63 downto 0);
      EMIOGPIOTN           : out std_logic_vector(63 downto 0);
      EMIOI2C0SCLO         : out std_ulogic;
      EMIOI2C0SCLTN        : out std_ulogic;
      EMIOI2C0SDAO         : out std_ulogic;
      EMIOI2C0SDATN        : out std_ulogic;
      EMIOI2C1SCLO         : out std_ulogic;
      EMIOI2C1SCLTN        : out std_ulogic;
      EMIOI2C1SDAO         : out std_ulogic;
      EMIOI2C1SDATN        : out std_ulogic;
      EMIOPJTAGTDO         : out std_ulogic;
      EMIOPJTAGTDTN        : out std_ulogic;
      EMIOSDIO0BUSPOW      : out std_ulogic;
      EMIOSDIO0BUSVOLT     : out std_logic_vector(2 downto 0);
      EMIOSDIO0CLK         : out std_ulogic;
      EMIOSDIO0CMDO        : out std_ulogic;
      EMIOSDIO0CMDTN       : out std_ulogic;
      EMIOSDIO0DATAO       : out std_logic_vector(3 downto 0);
      EMIOSDIO0DATATN      : out std_logic_vector(3 downto 0);
      EMIOSDIO0LED         : out std_ulogic;
      EMIOSDIO1BUSPOW      : out std_ulogic;
      EMIOSDIO1BUSVOLT     : out std_logic_vector(2 downto 0);
      EMIOSDIO1CLK         : out std_ulogic;
      EMIOSDIO1CMDO        : out std_ulogic;
      EMIOSDIO1CMDTN       : out std_ulogic;
      EMIOSDIO1DATAO       : out std_logic_vector(3 downto 0);
      EMIOSDIO1DATATN      : out std_logic_vector(3 downto 0);
      EMIOSDIO1LED         : out std_ulogic;
      EMIOSPI0MO           : out std_ulogic;
      EMIOSPI0MOTN         : out std_ulogic;
      EMIOSPI0SCLKO        : out std_ulogic;
      EMIOSPI0SCLKTN       : out std_ulogic;
      EMIOSPI0SO           : out std_ulogic;
      EMIOSPI0SSNTN        : out std_ulogic;
      EMIOSPI0SSON         : out std_logic_vector(2 downto 0);
      EMIOSPI0STN          : out std_ulogic;
      EMIOSPI1MO           : out std_ulogic;
      EMIOSPI1MOTN         : out std_ulogic;
      EMIOSPI1SCLKO        : out std_ulogic;
      EMIOSPI1SCLKTN       : out std_ulogic;
      EMIOSPI1SO           : out std_ulogic;
      EMIOSPI1SSNTN        : out std_ulogic;
      EMIOSPI1SSON         : out std_logic_vector(2 downto 0);
      EMIOSPI1STN          : out std_ulogic;
      EMIOTRACECTL         : out std_ulogic;
      EMIOTRACEDATA        : out std_logic_vector(31 downto 0);
      EMIOTTC0WAVEO        : out std_logic_vector(2 downto 0);
      EMIOTTC1WAVEO        : out std_logic_vector(2 downto 0);
      EMIOUART0DTRN        : out std_ulogic;
      EMIOUART0RTSN        : out std_ulogic;
      EMIOUART0TX          : out std_ulogic;
      EMIOUART1DTRN        : out std_ulogic;
      EMIOUART1RTSN        : out std_ulogic;
      EMIOUART1TX          : out std_ulogic;
      EMIOUSB0PORTINDCTL   : out std_logic_vector(1 downto 0);
      EMIOUSB0VBUSPWRSELECT : out std_ulogic;
      EMIOUSB1PORTINDCTL   : out std_logic_vector(1 downto 0);
      EMIOUSB1VBUSPWRSELECT : out std_ulogic;
      EMIOWDTRSTO          : out std_ulogic;
      EVENTEVENTO          : out std_ulogic;
      EVENTSTANDBYWFE      : out std_logic_vector(1 downto 0);
      EVENTSTANDBYWFI      : out std_logic_vector(1 downto 0);
      FCLKCLK              : out std_logic_vector(3 downto 0);
      FCLKRESETN           : out std_logic_vector(3 downto 0);
      FTMTF2PTRIGACK       : out std_logic_vector(3 downto 0);
      FTMTP2FDEBUG         : out std_logic_vector(31 downto 0);
      FTMTP2FTRIG          : out std_logic_vector(3 downto 0);
      IRQP2F               : out std_logic_vector(28 downto 0);
      MAXIGP0ARADDR        : out std_logic_vector(31 downto 0);
      MAXIGP0ARBURST       : out std_logic_vector(1 downto 0);
      MAXIGP0ARCACHE       : out std_logic_vector(3 downto 0);
      MAXIGP0ARESETN       : out std_ulogic;
      MAXIGP0ARID          : out std_logic_vector(11 downto 0);
      MAXIGP0ARLEN         : out std_logic_vector(3 downto 0);
      MAXIGP0ARLOCK        : out std_logic_vector(1 downto 0);
      MAXIGP0ARPROT        : out std_logic_vector(2 downto 0);
      MAXIGP0ARQOS         : out std_logic_vector(3 downto 0);
      MAXIGP0ARSIZE        : out std_logic_vector(1 downto 0);
      MAXIGP0ARVALID       : out std_ulogic;
      MAXIGP0AWADDR        : out std_logic_vector(31 downto 0);
      MAXIGP0AWBURST       : out std_logic_vector(1 downto 0);
      MAXIGP0AWCACHE       : out std_logic_vector(3 downto 0);
      MAXIGP0AWID          : out std_logic_vector(11 downto 0);
      MAXIGP0AWLEN         : out std_logic_vector(3 downto 0);
      MAXIGP0AWLOCK        : out std_logic_vector(1 downto 0);
      MAXIGP0AWPROT        : out std_logic_vector(2 downto 0);
      MAXIGP0AWQOS         : out std_logic_vector(3 downto 0);
      MAXIGP0AWSIZE        : out std_logic_vector(1 downto 0);
      MAXIGP0AWVALID       : out std_ulogic;
      MAXIGP0BREADY        : out std_ulogic;
      MAXIGP0RREADY        : out std_ulogic;
      MAXIGP0WDATA         : out std_logic_vector(31 downto 0);
      MAXIGP0WID           : out std_logic_vector(11 downto 0);
      MAXIGP0WLAST         : out std_ulogic;
      MAXIGP0WSTRB         : out std_logic_vector(3 downto 0);
      MAXIGP0WVALID        : out std_ulogic;
      MAXIGP1ARADDR        : out std_logic_vector(31 downto 0);
      MAXIGP1ARBURST       : out std_logic_vector(1 downto 0);
      MAXIGP1ARCACHE       : out std_logic_vector(3 downto 0);
      MAXIGP1ARESETN       : out std_ulogic;
      MAXIGP1ARID          : out std_logic_vector(11 downto 0);
      MAXIGP1ARLEN         : out std_logic_vector(3 downto 0);
      MAXIGP1ARLOCK        : out std_logic_vector(1 downto 0);
      MAXIGP1ARPROT        : out std_logic_vector(2 downto 0);
      MAXIGP1ARQOS         : out std_logic_vector(3 downto 0);
      MAXIGP1ARSIZE        : out std_logic_vector(1 downto 0);
      MAXIGP1ARVALID       : out std_ulogic;
      MAXIGP1AWADDR        : out std_logic_vector(31 downto 0);
      MAXIGP1AWBURST       : out std_logic_vector(1 downto 0);
      MAXIGP1AWCACHE       : out std_logic_vector(3 downto 0);
      MAXIGP1AWID          : out std_logic_vector(11 downto 0);
      MAXIGP1AWLEN         : out std_logic_vector(3 downto 0);
      MAXIGP1AWLOCK        : out std_logic_vector(1 downto 0);
      MAXIGP1AWPROT        : out std_logic_vector(2 downto 0);
      MAXIGP1AWQOS         : out std_logic_vector(3 downto 0);
      MAXIGP1AWSIZE        : out std_logic_vector(1 downto 0);
      MAXIGP1AWVALID       : out std_ulogic;
      MAXIGP1BREADY        : out std_ulogic;
      MAXIGP1RREADY        : out std_ulogic;
      MAXIGP1WDATA         : out std_logic_vector(31 downto 0);
      MAXIGP1WID           : out std_logic_vector(11 downto 0);
      MAXIGP1WLAST         : out std_ulogic;
      MAXIGP1WSTRB         : out std_logic_vector(3 downto 0);
      MAXIGP1WVALID        : out std_ulogic;
      SAXIACPARESETN       : out std_ulogic;
      SAXIACPARREADY       : out std_ulogic;
      SAXIACPAWREADY       : out std_ulogic;
      SAXIACPBID           : out std_logic_vector(2 downto 0);
      SAXIACPBRESP         : out std_logic_vector(1 downto 0);
      SAXIACPBVALID        : out std_ulogic;
      SAXIACPRDATA         : out std_logic_vector(63 downto 0);
      SAXIACPRID           : out std_logic_vector(2 downto 0);
      SAXIACPRLAST         : out std_ulogic;
      SAXIACPRRESP         : out std_logic_vector(1 downto 0);
      SAXIACPRVALID        : out std_ulogic;
      SAXIACPWREADY        : out std_ulogic;
      SAXIGP0ARESETN       : out std_ulogic;
      SAXIGP0ARREADY       : out std_ulogic;
      SAXIGP0AWREADY       : out std_ulogic;
      SAXIGP0BID           : out std_logic_vector(5 downto 0);
      SAXIGP0BRESP         : out std_logic_vector(1 downto 0);
      SAXIGP0BVALID        : out std_ulogic;
      SAXIGP0RDATA         : out std_logic_vector(31 downto 0);
      SAXIGP0RID           : out std_logic_vector(5 downto 0);
      SAXIGP0RLAST         : out std_ulogic;
      SAXIGP0RRESP         : out std_logic_vector(1 downto 0);
      SAXIGP0RVALID        : out std_ulogic;
      SAXIGP0WREADY        : out std_ulogic;
      SAXIGP1ARESETN       : out std_ulogic;
      SAXIGP1ARREADY       : out std_ulogic;
      SAXIGP1AWREADY       : out std_ulogic;
      SAXIGP1BID           : out std_logic_vector(5 downto 0);
      SAXIGP1BRESP         : out std_logic_vector(1 downto 0);
      SAXIGP1BVALID        : out std_ulogic;
      SAXIGP1RDATA         : out std_logic_vector(31 downto 0);
      SAXIGP1RID           : out std_logic_vector(5 downto 0);
      SAXIGP1RLAST         : out std_ulogic;
      SAXIGP1RRESP         : out std_logic_vector(1 downto 0);
      SAXIGP1RVALID        : out std_ulogic;
      SAXIGP1WREADY        : out std_ulogic;
      SAXIHP0ARESETN       : out std_ulogic;
      SAXIHP0ARREADY       : out std_ulogic;
      SAXIHP0AWREADY       : out std_ulogic;
      SAXIHP0BID           : out std_logic_vector(5 downto 0);
      SAXIHP0BRESP         : out std_logic_vector(1 downto 0);
      SAXIHP0BVALID        : out std_ulogic;
      SAXIHP0RACOUNT       : out std_logic_vector(2 downto 0);
      SAXIHP0RCOUNT        : out std_logic_vector(7 downto 0);
      SAXIHP0RDATA         : out std_logic_vector(63 downto 0);
      SAXIHP0RID           : out std_logic_vector(5 downto 0);
      SAXIHP0RLAST         : out std_ulogic;
      SAXIHP0RRESP         : out std_logic_vector(1 downto 0);
      SAXIHP0RVALID        : out std_ulogic;
      SAXIHP0WACOUNT       : out std_logic_vector(5 downto 0);
      SAXIHP0WCOUNT        : out std_logic_vector(7 downto 0);
      SAXIHP0WREADY        : out std_ulogic;
      SAXIHP1ARESETN       : out std_ulogic;
      SAXIHP1ARREADY       : out std_ulogic;
      SAXIHP1AWREADY       : out std_ulogic;
      SAXIHP1BID           : out std_logic_vector(5 downto 0);
      SAXIHP1BRESP         : out std_logic_vector(1 downto 0);
      SAXIHP1BVALID        : out std_ulogic;
      SAXIHP1RACOUNT       : out std_logic_vector(2 downto 0);
      SAXIHP1RCOUNT        : out std_logic_vector(7 downto 0);
      SAXIHP1RDATA         : out std_logic_vector(63 downto 0);
      SAXIHP1RID           : out std_logic_vector(5 downto 0);
      SAXIHP1RLAST         : out std_ulogic;
      SAXIHP1RRESP         : out std_logic_vector(1 downto 0);
      SAXIHP1RVALID        : out std_ulogic;
      SAXIHP1WACOUNT       : out std_logic_vector(5 downto 0);
      SAXIHP1WCOUNT        : out std_logic_vector(7 downto 0);
      SAXIHP1WREADY        : out std_ulogic;
      SAXIHP2ARESETN       : out std_ulogic;
      SAXIHP2ARREADY       : out std_ulogic;
      SAXIHP2AWREADY       : out std_ulogic;
      SAXIHP2BID           : out std_logic_vector(5 downto 0);
      SAXIHP2BRESP         : out std_logic_vector(1 downto 0);
      SAXIHP2BVALID        : out std_ulogic;
      SAXIHP2RACOUNT       : out std_logic_vector(2 downto 0);
      SAXIHP2RCOUNT        : out std_logic_vector(7 downto 0);
      SAXIHP2RDATA         : out std_logic_vector(63 downto 0);
      SAXIHP2RID           : out std_logic_vector(5 downto 0);
      SAXIHP2RLAST         : out std_ulogic;
      SAXIHP2RRESP         : out std_logic_vector(1 downto 0);
      SAXIHP2RVALID        : out std_ulogic;
      SAXIHP2WACOUNT       : out std_logic_vector(5 downto 0);
      SAXIHP2WCOUNT        : out std_logic_vector(7 downto 0);
      SAXIHP2WREADY        : out std_ulogic;
      SAXIHP3ARESETN       : out std_ulogic;
      SAXIHP3ARREADY       : out std_ulogic;
      SAXIHP3AWREADY       : out std_ulogic;
      SAXIHP3BID           : out std_logic_vector(5 downto 0);
      SAXIHP3BRESP         : out std_logic_vector(1 downto 0);
      SAXIHP3BVALID        : out std_ulogic;
      SAXIHP3RACOUNT       : out std_logic_vector(2 downto 0);
      SAXIHP3RCOUNT        : out std_logic_vector(7 downto 0);
      SAXIHP3RDATA         : out std_logic_vector(63 downto 0);
      SAXIHP3RID           : out std_logic_vector(5 downto 0);
      SAXIHP3RLAST         : out std_ulogic;
      SAXIHP3RRESP         : out std_logic_vector(1 downto 0);
      SAXIHP3RVALID        : out std_ulogic;
      SAXIHP3WACOUNT       : out std_logic_vector(5 downto 0);
      SAXIHP3WCOUNT        : out std_logic_vector(7 downto 0);
      SAXIHP3WREADY        : out std_ulogic;
      DDRA                 : inout std_logic_vector(14 downto 0);
      DDRBA                : inout std_logic_vector(2 downto 0);
      DDRCASB              : inout std_ulogic;
      DDRCKE               : inout std_ulogic;
      DDRCKN               : inout std_ulogic;
      DDRCKP               : inout std_ulogic;
      DDRCSB               : inout std_ulogic;
      DDRDM                : inout std_logic_vector(3 downto 0);
      DDRDQ                : inout std_logic_vector(31 downto 0);
      DDRDQSN              : inout std_logic_vector(3 downto 0);
      DDRDQSP              : inout std_logic_vector(3 downto 0);
      DDRDRSTB             : inout std_ulogic;
      DDRODT               : inout std_ulogic;
      DDRRASB              : inout std_ulogic;
      DDRVRN               : inout std_ulogic;
      DDRVRP               : inout std_ulogic;
      DDRWEB               : inout std_ulogic;
      MIO                  : inout std_logic_vector(53 downto 0);
      PSCLK                : inout std_ulogic;
      PSPORB               : inout std_ulogic;
      PSSRSTB              : inout std_ulogic;
      DDRARB               : in std_logic_vector(3 downto 0);
      DMA0ACLK             : in std_ulogic;
      DMA0DAREADY          : in std_ulogic;
      DMA0DRLAST           : in std_ulogic;
      DMA0DRTYPE           : in std_logic_vector(1 downto 0);
      DMA0DRVALID          : in std_ulogic;
      DMA1ACLK             : in std_ulogic;
      DMA1DAREADY          : in std_ulogic;
      DMA1DRLAST           : in std_ulogic;
      DMA1DRTYPE           : in std_logic_vector(1 downto 0);
      DMA1DRVALID          : in std_ulogic;
      DMA2ACLK             : in std_ulogic;
      DMA2DAREADY          : in std_ulogic;
      DMA2DRLAST           : in std_ulogic;
      DMA2DRTYPE           : in std_logic_vector(1 downto 0);
      DMA2DRVALID          : in std_ulogic;
      DMA3ACLK             : in std_ulogic;
      DMA3DAREADY          : in std_ulogic;
      DMA3DRLAST           : in std_ulogic;
      DMA3DRTYPE           : in std_logic_vector(1 downto 0);
      DMA3DRVALID          : in std_ulogic;
      EMIOCAN0PHYRX        : in std_ulogic;
      EMIOCAN1PHYRX        : in std_ulogic;
      EMIOENET0EXTINTIN    : in std_ulogic;
      EMIOENET0GMIICOL     : in std_ulogic;
      EMIOENET0GMIICRS     : in std_ulogic;
      EMIOENET0GMIIRXCLK   : in std_ulogic;
      EMIOENET0GMIIRXD     : in std_logic_vector(7 downto 0);
      EMIOENET0GMIIRXDV    : in std_ulogic;
      EMIOENET0GMIIRXER    : in std_ulogic;
      EMIOENET0GMIITXCLK   : in std_ulogic;
      EMIOENET0MDIOI       : in std_ulogic;
      EMIOENET1EXTINTIN    : in std_ulogic;
      EMIOENET1GMIICOL     : in std_ulogic;
      EMIOENET1GMIICRS     : in std_ulogic;
      EMIOENET1GMIIRXCLK   : in std_ulogic;
      EMIOENET1GMIIRXD     : in std_logic_vector(7 downto 0);
      EMIOENET1GMIIRXDV    : in std_ulogic;
      EMIOENET1GMIIRXER    : in std_ulogic;
      EMIOENET1GMIITXCLK   : in std_ulogic;
      EMIOENET1MDIOI       : in std_ulogic;
      EMIOGPIOI            : in std_logic_vector(63 downto 0);
      EMIOI2C0SCLI         : in std_ulogic;
      EMIOI2C0SDAI         : in std_ulogic;
      EMIOI2C1SCLI         : in std_ulogic;
      EMIOI2C1SDAI         : in std_ulogic;
      EMIOPJTAGTCK         : in std_ulogic;
      EMIOPJTAGTDI         : in std_ulogic;
      EMIOPJTAGTMS         : in std_ulogic;
      EMIOSDIO0CDN         : in std_ulogic;
      EMIOSDIO0CLKFB       : in std_ulogic;
      EMIOSDIO0CMDI        : in std_ulogic;
      EMIOSDIO0DATAI       : in std_logic_vector(3 downto 0);
      EMIOSDIO0WP          : in std_ulogic;
      EMIOSDIO1CDN         : in std_ulogic;
      EMIOSDIO1CLKFB       : in std_ulogic;
      EMIOSDIO1CMDI        : in std_ulogic;
      EMIOSDIO1DATAI       : in std_logic_vector(3 downto 0);
      EMIOSDIO1WP          : in std_ulogic;
      EMIOSPI0MI           : in std_ulogic;
      EMIOSPI0SCLKI        : in std_ulogic;
      EMIOSPI0SI           : in std_ulogic;
      EMIOSPI0SSIN         : in std_ulogic;
      EMIOSPI1MI           : in std_ulogic;
      EMIOSPI1SCLKI        : in std_ulogic;
      EMIOSPI1SI           : in std_ulogic;
      EMIOSPI1SSIN         : in std_ulogic;
      EMIOSRAMINTIN        : in std_ulogic;
      EMIOTRACECLK         : in std_ulogic;
      EMIOTTC0CLKI         : in std_logic_vector(2 downto 0);
      EMIOTTC1CLKI         : in std_logic_vector(2 downto 0);
      EMIOUART0CTSN        : in std_ulogic;
      EMIOUART0DCDN        : in std_ulogic;
      EMIOUART0DSRN        : in std_ulogic;
      EMIOUART0RIN         : in std_ulogic;
      EMIOUART0RX          : in std_ulogic;
      EMIOUART1CTSN        : in std_ulogic;
      EMIOUART1DCDN        : in std_ulogic;
      EMIOUART1DSRN        : in std_ulogic;
      EMIOUART1RIN         : in std_ulogic;
      EMIOUART1RX          : in std_ulogic;
      EMIOUSB0VBUSPWRFAULT : in std_ulogic;
      EMIOUSB1VBUSPWRFAULT : in std_ulogic;
      EMIOWDTCLKI          : in std_ulogic;
      EVENTEVENTI          : in std_ulogic;
      FCLKCLKTRIGN         : in std_logic_vector(3 downto 0);
      FPGAIDLEN            : in std_ulogic;
      FTMDTRACEINATID      : in std_logic_vector(3 downto 0);
      FTMDTRACEINCLOCK     : in std_ulogic;
      FTMDTRACEINDATA      : in std_logic_vector(31 downto 0);
      FTMDTRACEINVALID     : in std_ulogic;
      FTMTF2PDEBUG         : in std_logic_vector(31 downto 0);
      FTMTF2PTRIG          : in std_logic_vector(3 downto 0);
      FTMTP2FTRIGACK       : in std_logic_vector(3 downto 0);
      IRQF2P               : in std_logic_vector(19 downto 0);
      MAXIGP0ACLK          : in std_ulogic;
      MAXIGP0ARREADY       : in std_ulogic;
      MAXIGP0AWREADY       : in std_ulogic;
      MAXIGP0BID           : in std_logic_vector(11 downto 0);
      MAXIGP0BRESP         : in std_logic_vector(1 downto 0);
      MAXIGP0BVALID        : in std_ulogic;
      MAXIGP0RDATA         : in std_logic_vector(31 downto 0);
      MAXIGP0RID           : in std_logic_vector(11 downto 0);
      MAXIGP0RLAST         : in std_ulogic;
      MAXIGP0RRESP         : in std_logic_vector(1 downto 0);
      MAXIGP0RVALID        : in std_ulogic;
      MAXIGP0WREADY        : in std_ulogic;
      MAXIGP1ACLK          : in std_ulogic;
      MAXIGP1ARREADY       : in std_ulogic;
      MAXIGP1AWREADY       : in std_ulogic;
      MAXIGP1BID           : in std_logic_vector(11 downto 0);
      MAXIGP1BRESP         : in std_logic_vector(1 downto 0);
      MAXIGP1BVALID        : in std_ulogic;
      MAXIGP1RDATA         : in std_logic_vector(31 downto 0);
      MAXIGP1RID           : in std_logic_vector(11 downto 0);
      MAXIGP1RLAST         : in std_ulogic;
      MAXIGP1RRESP         : in std_logic_vector(1 downto 0);
      MAXIGP1RVALID        : in std_ulogic;
      MAXIGP1WREADY        : in std_ulogic;
      SAXIACPACLK          : in std_ulogic;
      SAXIACPARADDR        : in std_logic_vector(31 downto 0);
      SAXIACPARBURST       : in std_logic_vector(1 downto 0);
      SAXIACPARCACHE       : in std_logic_vector(3 downto 0);
      SAXIACPARID          : in std_logic_vector(2 downto 0);
      SAXIACPARLEN         : in std_logic_vector(3 downto 0);
      SAXIACPARLOCK        : in std_logic_vector(1 downto 0);
      SAXIACPARPROT        : in std_logic_vector(2 downto 0);
      SAXIACPARQOS         : in std_logic_vector(3 downto 0);
      SAXIACPARSIZE        : in std_logic_vector(1 downto 0);
      SAXIACPARUSER        : in std_logic_vector(4 downto 0);
      SAXIACPARVALID       : in std_ulogic;
      SAXIACPAWADDR        : in std_logic_vector(31 downto 0);
      SAXIACPAWBURST       : in std_logic_vector(1 downto 0);
      SAXIACPAWCACHE       : in std_logic_vector(3 downto 0);
      SAXIACPAWID          : in std_logic_vector(2 downto 0);
      SAXIACPAWLEN         : in std_logic_vector(3 downto 0);
      SAXIACPAWLOCK        : in std_logic_vector(1 downto 0);
      SAXIACPAWPROT        : in std_logic_vector(2 downto 0);
      SAXIACPAWQOS         : in std_logic_vector(3 downto 0);
      SAXIACPAWSIZE        : in std_logic_vector(1 downto 0);
      SAXIACPAWUSER        : in std_logic_vector(4 downto 0);
      SAXIACPAWVALID       : in std_ulogic;
      SAXIACPBREADY        : in std_ulogic;
      SAXIACPRREADY        : in std_ulogic;
      SAXIACPWDATA         : in std_logic_vector(63 downto 0);
      SAXIACPWID           : in std_logic_vector(2 downto 0);
      SAXIACPWLAST         : in std_ulogic;
      SAXIACPWSTRB         : in std_logic_vector(7 downto 0);
      SAXIACPWVALID        : in std_ulogic;
      SAXIGP0ACLK          : in std_ulogic;
      SAXIGP0ARADDR        : in std_logic_vector(31 downto 0);
      SAXIGP0ARBURST       : in std_logic_vector(1 downto 0);
      SAXIGP0ARCACHE       : in std_logic_vector(3 downto 0);
      SAXIGP0ARID          : in std_logic_vector(5 downto 0);
      SAXIGP0ARLEN         : in std_logic_vector(3 downto 0);
      SAXIGP0ARLOCK        : in std_logic_vector(1 downto 0);
      SAXIGP0ARPROT        : in std_logic_vector(2 downto 0);
      SAXIGP0ARQOS         : in std_logic_vector(3 downto 0);
      SAXIGP0ARSIZE        : in std_logic_vector(1 downto 0);
      SAXIGP0ARVALID       : in std_ulogic;
      SAXIGP0AWADDR        : in std_logic_vector(31 downto 0);
      SAXIGP0AWBURST       : in std_logic_vector(1 downto 0);
      SAXIGP0AWCACHE       : in std_logic_vector(3 downto 0);
      SAXIGP0AWID          : in std_logic_vector(5 downto 0);
      SAXIGP0AWLEN         : in std_logic_vector(3 downto 0);
      SAXIGP0AWLOCK        : in std_logic_vector(1 downto 0);
      SAXIGP0AWPROT        : in std_logic_vector(2 downto 0);
      SAXIGP0AWQOS         : in std_logic_vector(3 downto 0);
      SAXIGP0AWSIZE        : in std_logic_vector(1 downto 0);
      SAXIGP0AWVALID       : in std_ulogic;
      SAXIGP0BREADY        : in std_ulogic;
      SAXIGP0RREADY        : in std_ulogic;
      SAXIGP0WDATA         : in std_logic_vector(31 downto 0);
      SAXIGP0WID           : in std_logic_vector(5 downto 0);
      SAXIGP0WLAST         : in std_ulogic;
      SAXIGP0WSTRB         : in std_logic_vector(3 downto 0);
      SAXIGP0WVALID        : in std_ulogic;
      SAXIGP1ACLK          : in std_ulogic;
      SAXIGP1ARADDR        : in std_logic_vector(31 downto 0);
      SAXIGP1ARBURST       : in std_logic_vector(1 downto 0);
      SAXIGP1ARCACHE       : in std_logic_vector(3 downto 0);
      SAXIGP1ARID          : in std_logic_vector(5 downto 0);
      SAXIGP1ARLEN         : in std_logic_vector(3 downto 0);
      SAXIGP1ARLOCK        : in std_logic_vector(1 downto 0);
      SAXIGP1ARPROT        : in std_logic_vector(2 downto 0);
      SAXIGP1ARQOS         : in std_logic_vector(3 downto 0);
      SAXIGP1ARSIZE        : in std_logic_vector(1 downto 0);
      SAXIGP1ARVALID       : in std_ulogic;
      SAXIGP1AWADDR        : in std_logic_vector(31 downto 0);
      SAXIGP1AWBURST       : in std_logic_vector(1 downto 0);
      SAXIGP1AWCACHE       : in std_logic_vector(3 downto 0);
      SAXIGP1AWID          : in std_logic_vector(5 downto 0);
      SAXIGP1AWLEN         : in std_logic_vector(3 downto 0);
      SAXIGP1AWLOCK        : in std_logic_vector(1 downto 0);
      SAXIGP1AWPROT        : in std_logic_vector(2 downto 0);
      SAXIGP1AWQOS         : in std_logic_vector(3 downto 0);
      SAXIGP1AWSIZE        : in std_logic_vector(1 downto 0);
      SAXIGP1AWVALID       : in std_ulogic;
      SAXIGP1BREADY        : in std_ulogic;
      SAXIGP1RREADY        : in std_ulogic;
      SAXIGP1WDATA         : in std_logic_vector(31 downto 0);
      SAXIGP1WID           : in std_logic_vector(5 downto 0);
      SAXIGP1WLAST         : in std_ulogic;
      SAXIGP1WSTRB         : in std_logic_vector(3 downto 0);
      SAXIGP1WVALID        : in std_ulogic;
      SAXIHP0ACLK          : in std_ulogic;
      SAXIHP0ARADDR        : in std_logic_vector(31 downto 0);
      SAXIHP0ARBURST       : in std_logic_vector(1 downto 0);
      SAXIHP0ARCACHE       : in std_logic_vector(3 downto 0);
      SAXIHP0ARID          : in std_logic_vector(5 downto 0);
      SAXIHP0ARLEN         : in std_logic_vector(3 downto 0);
      SAXIHP0ARLOCK        : in std_logic_vector(1 downto 0);
      SAXIHP0ARPROT        : in std_logic_vector(2 downto 0);
      SAXIHP0ARQOS         : in std_logic_vector(3 downto 0);
      SAXIHP0ARSIZE        : in std_logic_vector(1 downto 0);
      SAXIHP0ARVALID       : in std_ulogic;
      SAXIHP0AWADDR        : in std_logic_vector(31 downto 0);
      SAXIHP0AWBURST       : in std_logic_vector(1 downto 0);
      SAXIHP0AWCACHE       : in std_logic_vector(3 downto 0);
      SAXIHP0AWID          : in std_logic_vector(5 downto 0);
      SAXIHP0AWLEN         : in std_logic_vector(3 downto 0);
      SAXIHP0AWLOCK        : in std_logic_vector(1 downto 0);
      SAXIHP0AWPROT        : in std_logic_vector(2 downto 0);
      SAXIHP0AWQOS         : in std_logic_vector(3 downto 0);
      SAXIHP0AWSIZE        : in std_logic_vector(1 downto 0);
      SAXIHP0AWVALID       : in std_ulogic;
      SAXIHP0BREADY        : in std_ulogic;
      SAXIHP0RDISSUECAP1EN : in std_ulogic;
      SAXIHP0RREADY        : in std_ulogic;
      SAXIHP0WDATA         : in std_logic_vector(63 downto 0);
      SAXIHP0WID           : in std_logic_vector(5 downto 0);
      SAXIHP0WLAST         : in std_ulogic;
      SAXIHP0WRISSUECAP1EN : in std_ulogic;
      SAXIHP0WSTRB         : in std_logic_vector(7 downto 0);
      SAXIHP0WVALID        : in std_ulogic;
      SAXIHP1ACLK          : in std_ulogic;
      SAXIHP1ARADDR        : in std_logic_vector(31 downto 0);
      SAXIHP1ARBURST       : in std_logic_vector(1 downto 0);
      SAXIHP1ARCACHE       : in std_logic_vector(3 downto 0);
      SAXIHP1ARID          : in std_logic_vector(5 downto 0);
      SAXIHP1ARLEN         : in std_logic_vector(3 downto 0);
      SAXIHP1ARLOCK        : in std_logic_vector(1 downto 0);
      SAXIHP1ARPROT        : in std_logic_vector(2 downto 0);
      SAXIHP1ARQOS         : in std_logic_vector(3 downto 0);
      SAXIHP1ARSIZE        : in std_logic_vector(1 downto 0);
      SAXIHP1ARVALID       : in std_ulogic;
      SAXIHP1AWADDR        : in std_logic_vector(31 downto 0);
      SAXIHP1AWBURST       : in std_logic_vector(1 downto 0);
      SAXIHP1AWCACHE       : in std_logic_vector(3 downto 0);
      SAXIHP1AWID          : in std_logic_vector(5 downto 0);
      SAXIHP1AWLEN         : in std_logic_vector(3 downto 0);
      SAXIHP1AWLOCK        : in std_logic_vector(1 downto 0);
      SAXIHP1AWPROT        : in std_logic_vector(2 downto 0);
      SAXIHP1AWQOS         : in std_logic_vector(3 downto 0);
      SAXIHP1AWSIZE        : in std_logic_vector(1 downto 0);
      SAXIHP1AWVALID       : in std_ulogic;
      SAXIHP1BREADY        : in std_ulogic;
      SAXIHP1RDISSUECAP1EN : in std_ulogic;
      SAXIHP1RREADY        : in std_ulogic;
      SAXIHP1WDATA         : in std_logic_vector(63 downto 0);
      SAXIHP1WID           : in std_logic_vector(5 downto 0);
      SAXIHP1WLAST         : in std_ulogic;
      SAXIHP1WRISSUECAP1EN : in std_ulogic;
      SAXIHP1WSTRB         : in std_logic_vector(7 downto 0);
      SAXIHP1WVALID        : in std_ulogic;
      SAXIHP2ACLK          : in std_ulogic;
      SAXIHP2ARADDR        : in std_logic_vector(31 downto 0);
      SAXIHP2ARBURST       : in std_logic_vector(1 downto 0);
      SAXIHP2ARCACHE       : in std_logic_vector(3 downto 0);
      SAXIHP2ARID          : in std_logic_vector(5 downto 0);
      SAXIHP2ARLEN         : in std_logic_vector(3 downto 0);
      SAXIHP2ARLOCK        : in std_logic_vector(1 downto 0);
      SAXIHP2ARPROT        : in std_logic_vector(2 downto 0);
      SAXIHP2ARQOS         : in std_logic_vector(3 downto 0);
      SAXIHP2ARSIZE        : in std_logic_vector(1 downto 0);
      SAXIHP2ARVALID       : in std_ulogic;
      SAXIHP2AWADDR        : in std_logic_vector(31 downto 0);
      SAXIHP2AWBURST       : in std_logic_vector(1 downto 0);
      SAXIHP2AWCACHE       : in std_logic_vector(3 downto 0);
      SAXIHP2AWID          : in std_logic_vector(5 downto 0);
      SAXIHP2AWLEN         : in std_logic_vector(3 downto 0);
      SAXIHP2AWLOCK        : in std_logic_vector(1 downto 0);
      SAXIHP2AWPROT        : in std_logic_vector(2 downto 0);
      SAXIHP2AWQOS         : in std_logic_vector(3 downto 0);
      SAXIHP2AWSIZE        : in std_logic_vector(1 downto 0);
      SAXIHP2AWVALID       : in std_ulogic;
      SAXIHP2BREADY        : in std_ulogic;
      SAXIHP2RDISSUECAP1EN : in std_ulogic;
      SAXIHP2RREADY        : in std_ulogic;
      SAXIHP2WDATA         : in std_logic_vector(63 downto 0);
      SAXIHP2WID           : in std_logic_vector(5 downto 0);
      SAXIHP2WLAST         : in std_ulogic;
      SAXIHP2WRISSUECAP1EN : in std_ulogic;
      SAXIHP2WSTRB         : in std_logic_vector(7 downto 0);
      SAXIHP2WVALID        : in std_ulogic;
      SAXIHP3ACLK          : in std_ulogic;
      SAXIHP3ARADDR        : in std_logic_vector(31 downto 0);
      SAXIHP3ARBURST       : in std_logic_vector(1 downto 0);
      SAXIHP3ARCACHE       : in std_logic_vector(3 downto 0);
      SAXIHP3ARID          : in std_logic_vector(5 downto 0);
      SAXIHP3ARLEN         : in std_logic_vector(3 downto 0);
      SAXIHP3ARLOCK        : in std_logic_vector(1 downto 0);
      SAXIHP3ARPROT        : in std_logic_vector(2 downto 0);
      SAXIHP3ARQOS         : in std_logic_vector(3 downto 0);
      SAXIHP3ARSIZE        : in std_logic_vector(1 downto 0);
      SAXIHP3ARVALID       : in std_ulogic;
      SAXIHP3AWADDR        : in std_logic_vector(31 downto 0);
      SAXIHP3AWBURST       : in std_logic_vector(1 downto 0);
      SAXIHP3AWCACHE       : in std_logic_vector(3 downto 0);
      SAXIHP3AWID          : in std_logic_vector(5 downto 0);
      SAXIHP3AWLEN         : in std_logic_vector(3 downto 0);
      SAXIHP3AWLOCK        : in std_logic_vector(1 downto 0);
      SAXIHP3AWPROT        : in std_logic_vector(2 downto 0);
      SAXIHP3AWQOS         : in std_logic_vector(3 downto 0);
      SAXIHP3AWSIZE        : in std_logic_vector(1 downto 0);
      SAXIHP3AWVALID       : in std_ulogic;
      SAXIHP3BREADY        : in std_ulogic;
      SAXIHP3RDISSUECAP1EN : in std_ulogic;
      SAXIHP3RREADY        : in std_ulogic;
      SAXIHP3WDATA         : in std_logic_vector(63 downto 0);
      SAXIHP3WID           : in std_logic_vector(5 downto 0);
      SAXIHP3WLAST         : in std_ulogic;
      SAXIHP3WRISSUECAP1EN : in std_ulogic;
      SAXIHP3WSTRB         : in std_logic_vector(7 downto 0);
      SAXIHP3WVALID        : in std_ulogic      
    );
  end PS7;

  architecture PS7_V of PS7 is
  
  begin
    process
      variable Message : line;
    begin
       Write ( Message, string'( "Warning on instance " ));
       Write ( Message, string'( PS7'INSTANCE_NAME));
       Write ( Message, string'(" The Zynq-7000 All Programmable SoC does not have a simulation model. Behavioral simulation of Zynq-7000 (e.g. Zynq PS7 block) is not supported in any simulator. Please use the AXI BFM simulation model to verify the AXI transactions" ));
       report Message.all;
       DEALLOCATE (Message);
    wait;   
    end process;
  end PS7_V;
